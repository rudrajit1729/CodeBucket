module Binary2Exs3(a,b);
input [3:0]a;
output [3:0]b;
assign b=a+3;
endmodule

